.include xor.spice
.include xor_high.spice
.include xor_multifinger.spice

Vs vdd gnd 2.5
VA A gnd 0 PULSE(0 2.5 14u 10n 10n 27u 56u 0)
VB B gnd 0 PULSE(0 2.5 15u 10n 10n 10u 20u 0)
X1 fxor_multi A B vdd XOR_MULTI
X2 fxor_low A B vdd XOR_LOW
X3 fxor_high A B vdd XOR_HIGH
.tran 1u 100u

.control
	run
	plot A, B
	plot fxor_multi, fxor_low, fxor_high
.endc
.end
