* SPICE3 file created from /home/nikoszaza/Desktop/VLSI/project/part1/dff_multifinger.ext - technology: scmos

.include 0.25_models.txt

.subckt DFF_MULTI Q Qbar D CLK Vdd
M1000 Qbar CLK a_30_n13# w_101_5# CMOSN w=4u l=2u
+  ad=92p pd=80u as=144p ps=96u
M1001 Gnd Qbar Q Gnd CMOSN w=8u l=2u
+  ad=324p pd=232u as=96p ps=56u
M1002 Vdd Q Qbar Vdd CMOSP w=6u l=2u
+  ad=792p pd=384u as=216p ps=120u
M1003 a_30_n13# DG Vdd Vdd CMOSP w=24u l=2u
+  ad=432p pd=192u as=0p ps=0u
M1004 DG CLK D Vdd CMOSP w=12u l=2u
+  ad=216p pd=120u as=144p ps=72u
M1005 Gnd a_30_n13# DG Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=92p ps=80u
M1006 DG CLKN D Gnd CMOSN w=4u l=2u
+  ad=0p pd=0u as=48p ps=40u
M1007 CLKN CLK Gnd Gnd CMOSN w=3u l=2u
+  ad=44p pd=40u as=0p ps=0u
M1008 Q Qbar Gnd Gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_30_n13# CLK Qbar w_101_5# CMOSN w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1010 Qbar Q Vdd Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1011 Vdd CLK CLKN Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=72p ps=48u
M1012 Vdd a_30_n13# DG Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1013 Gnd Q Qbar Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_30_n13# DG Gnd Gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q Qbar Vdd Vdd CMOSP w=24u l=2u
+  ad=288p pd=120u as=0p ps=0u
M1016 Gnd a_30_n13# DG Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1017 Qbar CLKN a_30_n13# w_99_n20# CMOSP w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1018 CLKN CLK Gnd Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1019 Qbar CLK a_30_n13# w_101_5# CMOSN w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1020 D CLKN DG Gnd CMOSN w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1021 DG a_30_n13# Vdd Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1022 Gnd DG a_30_n13# Gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_30_n13# DG Vdd Vdd CMOSP w=24u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1024 Vdd Qbar Q Vdd CMOSP w=24u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1025 DG CLKN D Gnd CMOSN w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_30_n13# CLKN Qbar w_99_n20# CMOSP w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1027 CLKN CLK Vdd Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_30_n13# DG Gnd Gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1029 DG CLK D Vdd CMOSP w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1030 Vdd a_30_n13# DG Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1031 Qbar Q Vdd Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1032 DG a_30_n13# Gnd Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1033 Vdd DG a_30_n13# Vdd CMOSP w=24u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q Qbar Gnd Gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1035 Gnd CLK CLKN Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1036 D CLK DG Vdd CMOSP w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q Qbar Vdd Vdd CMOSP w=24u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1038 Qbar CLKN a_30_n13# w_99_n20# CMOSP w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1039 CLKN CLK Vdd Vdd CMOSP w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1040 Qbar Q Gnd Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1041 Qbar Q Gnd Gnd CMOSN w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 a_30_n13# Vdd 17.95fF
C1 Qbar Vdd 7.13fF
C2 w_101_5# Qbar 3.01fF
C3 CLKN DG 2.16fF
C4 CLKN w_99_n20# 4.36fF
C5 CLK Gnd 7.47fF
C6 Q Gnd 6.75fF
C7 CLKN Gnd 51.16fF
C8 Gnd DG 24.60fF
C9 CLK Vdd 63.73fF
C10 Q Vdd 6.75fF
C11 Gnd a_30_n13# 8.56fF
C12 Qbar Gnd 21.01fF
C13 CLK w_101_5# 6.83fF
C14 DG Vdd 11.84fF
C15 Q 0 16.11fF
C16 Qbar 0 23.91fF
C17 a_30_n13# 0 22.96fF
.ends DFF_MULTI
