* SPICE3 file created from /home/nikoszaza/Desktop/VLSI/project/xnor.ext - technology: scmos

.include 0.25_models.txt

.subckt XNOR_LOW xnor A B vdd
M1000 a_1_n3# a_n31_n33# xnor vdd CMOSP w=20u l=2u
+  ad=340p pd=114u as=120p ps=52u
M1001 a_n31_n33# A gnd gnd CMOSN w=4u l=2u
+  ad=24p pd=20u as=136p ps=78u
M1002 a_n7_n33# B xnor gnd CMOSN w=8u l=2u
+  ad=72p pd=34u as=152p ps=70u
M1003 gnd a_n31_n33# a_n7_n33# gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 gnd B a_29_n42# gnd CMOSN w=4u l=2u
+  ad=0p pd=0u as=24p ps=20u
M1005 vdd A a_n17_n3# vdd CMOSP w=20u l=2u
+  ad=240p pd=116u as=300p ps=110u
M1006 xnor a_29_n42# a_17_n33# gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=96p ps=40u
M1007 vdd B a_29_n42# vdd CMOSP w=10u l=2u
+  ad=0p pd=0u as=60p ps=32u
M1008 a_17_n33# A gnd gnd CMOSN w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_n31_n33# A vdd vdd CMOSP w=10u l=2u
+  ad=60p pd=32u as=0p ps=0u
M1010 a_1_n3# a_29_n42# vdd vdd CMOSP w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1011 xnor B a_n17_n3# vdd CMOSP w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 vdd B 4.53fF
C1 gnd B 28.25fF
C2 a_1_n3# a_n17_n3# 3.76fF
C3 a_1_n3# vdd 3.29fF
C4 vdd a_29_n42# 2.84fF
C5 vdd A 22.06fF
C6 vdd a_n31_n33# 15.41fF
C7 gnd xnor 5.55fF
C8 gnd a_29_n42# 17.01fF
C9 gnd A 9.05fF
C10 gnd a_n31_n33# 6.68fF
C11 xnor 0 4.79fF
C12 a_29_n42# 0 6.43fF
C13 a_n31_n33# 0 6.80fF
.ends XNOR_LOW
