.include /home/znikolaos-g/VLSI/Project/Part2/dff.spice
.include dff_high.spice
.include dff_multifinger.spice

Vs vdd gnd 2.5
Vin D gnd 0 PULSE(0 2.5 14u 10n 10n 27u 56u 0)
Vclk clk gnd 0 PULSE(0 2.5 15u 10n 10n 10u 20u 0)
X1 Q_multi Qbar_multi D CLK vdd DFF_MULTI
X2 Q_high Qbar_high D CLK vdd DFF_HIGH
X3 Q_low Qbar_low D CLK vdd DFF_LOW

.tran 1u 100u 
.control
	run
	plot v(Q_low), v(D), v(Q_high), v(Q_multi)
	plot v(clk), v(D)
.endc
.end
